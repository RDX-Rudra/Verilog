mudule dlatch (output reg Q, Qn,
    input c, d
);
    
endmodule